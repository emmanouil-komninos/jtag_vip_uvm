`include "jtag_sequence_item.svh"
`include "jtag_config.svh"

`include "jtag_sequence_lib.svh"

`include "jtag_sequencer.svh"
`include "jtag_driver.svh"
`include "jtag_agent.svh"

`include "jtag_env.svh"
